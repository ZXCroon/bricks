library verilog;
use verilog.vl_types.all;
entity ball_move_computation is
    port(
        clk             : in     vl_logic;
        \ball.position_1_0\: in     vl_logic;
        \ball.position_1_1\: in     vl_logic;
        \ball.position_1_2\: in     vl_logic;
        \ball.position_1_3\: in     vl_logic;
        \ball.position_1_4\: in     vl_logic;
        \ball.position_1_5\: in     vl_logic;
        \ball.position_1_6\: in     vl_logic;
        \ball.position_1_7\: in     vl_logic;
        \ball.position_1_8\: in     vl_logic;
        \ball.position_1_9\: in     vl_logic;
        \ball.position_1_10\: in     vl_logic;
        \ball.position_1_11\: in     vl_logic;
        \ball.position_1_12\: in     vl_logic;
        \ball.position_1_13\: in     vl_logic;
        \ball.position_1_14\: in     vl_logic;
        \ball.position_1_15\: in     vl_logic;
        \ball.position_1_16\: in     vl_logic;
        \ball.position_1_17\: in     vl_logic;
        \ball.position_1_18\: in     vl_logic;
        \ball.position_1_19\: in     vl_logic;
        \ball.position_1_20\: in     vl_logic;
        \ball.position_1_21\: in     vl_logic;
        \ball.position_1_22\: in     vl_logic;
        \ball.position_1_23\: in     vl_logic;
        \ball.position_1_24\: in     vl_logic;
        \ball.position_1_25\: in     vl_logic;
        \ball.position_1_26\: in     vl_logic;
        \ball.position_1_27\: in     vl_logic;
        \ball.position_1_28\: in     vl_logic;
        \ball.position_1_29\: in     vl_logic;
        \ball.position_1_30\: in     vl_logic;
        \ball.position_1_31\: in     vl_logic;
        \ball.position_0_0\: in     vl_logic;
        \ball.position_0_1\: in     vl_logic;
        \ball.position_0_2\: in     vl_logic;
        \ball.position_0_3\: in     vl_logic;
        \ball.position_0_4\: in     vl_logic;
        \ball.position_0_5\: in     vl_logic;
        \ball.position_0_6\: in     vl_logic;
        \ball.position_0_7\: in     vl_logic;
        \ball.position_0_8\: in     vl_logic;
        \ball.position_0_9\: in     vl_logic;
        \ball.position_0_10\: in     vl_logic;
        \ball.position_0_11\: in     vl_logic;
        \ball.position_0_12\: in     vl_logic;
        \ball.position_0_13\: in     vl_logic;
        \ball.position_0_14\: in     vl_logic;
        \ball.position_0_15\: in     vl_logic;
        \ball.position_0_16\: in     vl_logic;
        \ball.position_0_17\: in     vl_logic;
        \ball.position_0_18\: in     vl_logic;
        \ball.position_0_19\: in     vl_logic;
        \ball.position_0_20\: in     vl_logic;
        \ball.position_0_21\: in     vl_logic;
        \ball.position_0_22\: in     vl_logic;
        \ball.position_0_23\: in     vl_logic;
        \ball.position_0_24\: in     vl_logic;
        \ball.position_0_25\: in     vl_logic;
        \ball.position_0_26\: in     vl_logic;
        \ball.position_0_27\: in     vl_logic;
        \ball.position_0_28\: in     vl_logic;
        \ball.position_0_29\: in     vl_logic;
        \ball.position_0_30\: in     vl_logic;
        \ball.position_0_31\: in     vl_logic;
        \ball.radius\   : in     vl_logic_vector(31 downto 0);
        velocity_1_31   : in     vl_logic;
        velocity_1_30   : in     vl_logic;
        velocity_1_29   : in     vl_logic;
        velocity_1_28   : in     vl_logic;
        velocity_1_27   : in     vl_logic;
        velocity_1_26   : in     vl_logic;
        velocity_1_25   : in     vl_logic;
        velocity_1_24   : in     vl_logic;
        velocity_1_23   : in     vl_logic;
        velocity_1_22   : in     vl_logic;
        velocity_1_21   : in     vl_logic;
        velocity_1_20   : in     vl_logic;
        velocity_1_19   : in     vl_logic;
        velocity_1_18   : in     vl_logic;
        velocity_1_17   : in     vl_logic;
        velocity_1_16   : in     vl_logic;
        velocity_1_15   : in     vl_logic;
        velocity_1_14   : in     vl_logic;
        velocity_1_13   : in     vl_logic;
        velocity_1_12   : in     vl_logic;
        velocity_1_11   : in     vl_logic;
        velocity_1_10   : in     vl_logic;
        velocity_1_9    : in     vl_logic;
        velocity_1_8    : in     vl_logic;
        velocity_1_7    : in     vl_logic;
        velocity_1_6    : in     vl_logic;
        velocity_1_5    : in     vl_logic;
        velocity_1_4    : in     vl_logic;
        velocity_1_3    : in     vl_logic;
        velocity_1_2    : in     vl_logic;
        velocity_1_1    : in     vl_logic;
        velocity_1_0    : in     vl_logic;
        velocity_0_31   : in     vl_logic;
        velocity_0_30   : in     vl_logic;
        velocity_0_29   : in     vl_logic;
        velocity_0_28   : in     vl_logic;
        velocity_0_27   : in     vl_logic;
        velocity_0_26   : in     vl_logic;
        velocity_0_25   : in     vl_logic;
        velocity_0_24   : in     vl_logic;
        velocity_0_23   : in     vl_logic;
        velocity_0_22   : in     vl_logic;
        velocity_0_21   : in     vl_logic;
        velocity_0_20   : in     vl_logic;
        velocity_0_19   : in     vl_logic;
        velocity_0_18   : in     vl_logic;
        velocity_0_17   : in     vl_logic;
        velocity_0_16   : in     vl_logic;
        velocity_0_15   : in     vl_logic;
        velocity_0_14   : in     vl_logic;
        velocity_0_13   : in     vl_logic;
        velocity_0_12   : in     vl_logic;
        velocity_0_11   : in     vl_logic;
        velocity_0_10   : in     vl_logic;
        velocity_0_9    : in     vl_logic;
        velocity_0_8    : in     vl_logic;
        velocity_0_7    : in     vl_logic;
        velocity_0_6    : in     vl_logic;
        velocity_0_5    : in     vl_logic;
        velocity_0_4    : in     vl_logic;
        velocity_0_3    : in     vl_logic;
        velocity_0_2    : in     vl_logic;
        velocity_0_1    : in     vl_logic;
        velocity_0_0    : in     vl_logic;
        \ball_next.position_1_0\: out    vl_logic;
        \ball_next.position_1_1\: out    vl_logic;
        \ball_next.position_1_2\: out    vl_logic;
        \ball_next.position_1_3\: out    vl_logic;
        \ball_next.position_1_4\: out    vl_logic;
        \ball_next.position_1_5\: out    vl_logic;
        \ball_next.position_1_6\: out    vl_logic;
        \ball_next.position_1_7\: out    vl_logic;
        \ball_next.position_1_8\: out    vl_logic;
        \ball_next.position_1_9\: out    vl_logic;
        \ball_next.position_1_10\: out    vl_logic;
        \ball_next.position_1_11\: out    vl_logic;
        \ball_next.position_1_12\: out    vl_logic;
        \ball_next.position_1_13\: out    vl_logic;
        \ball_next.position_1_14\: out    vl_logic;
        \ball_next.position_1_15\: out    vl_logic;
        \ball_next.position_1_16\: out    vl_logic;
        \ball_next.position_1_17\: out    vl_logic;
        \ball_next.position_1_18\: out    vl_logic;
        \ball_next.position_1_19\: out    vl_logic;
        \ball_next.position_1_20\: out    vl_logic;
        \ball_next.position_1_21\: out    vl_logic;
        \ball_next.position_1_22\: out    vl_logic;
        \ball_next.position_1_23\: out    vl_logic;
        \ball_next.position_1_24\: out    vl_logic;
        \ball_next.position_1_25\: out    vl_logic;
        \ball_next.position_1_26\: out    vl_logic;
        \ball_next.position_1_27\: out    vl_logic;
        \ball_next.position_1_28\: out    vl_logic;
        \ball_next.position_1_29\: out    vl_logic;
        \ball_next.position_1_30\: out    vl_logic;
        \ball_next.position_1_31\: out    vl_logic;
        \ball_next.position_0_0\: out    vl_logic;
        \ball_next.position_0_1\: out    vl_logic;
        \ball_next.position_0_2\: out    vl_logic;
        \ball_next.position_0_3\: out    vl_logic;
        \ball_next.position_0_4\: out    vl_logic;
        \ball_next.position_0_5\: out    vl_logic;
        \ball_next.position_0_6\: out    vl_logic;
        \ball_next.position_0_7\: out    vl_logic;
        \ball_next.position_0_8\: out    vl_logic;
        \ball_next.position_0_9\: out    vl_logic;
        \ball_next.position_0_10\: out    vl_logic;
        \ball_next.position_0_11\: out    vl_logic;
        \ball_next.position_0_12\: out    vl_logic;
        \ball_next.position_0_13\: out    vl_logic;
        \ball_next.position_0_14\: out    vl_logic;
        \ball_next.position_0_15\: out    vl_logic;
        \ball_next.position_0_16\: out    vl_logic;
        \ball_next.position_0_17\: out    vl_logic;
        \ball_next.position_0_18\: out    vl_logic;
        \ball_next.position_0_19\: out    vl_logic;
        \ball_next.position_0_20\: out    vl_logic;
        \ball_next.position_0_21\: out    vl_logic;
        \ball_next.position_0_22\: out    vl_logic;
        \ball_next.position_0_23\: out    vl_logic;
        \ball_next.position_0_24\: out    vl_logic;
        \ball_next.position_0_25\: out    vl_logic;
        \ball_next.position_0_26\: out    vl_logic;
        \ball_next.position_0_27\: out    vl_logic;
        \ball_next.position_0_28\: out    vl_logic;
        \ball_next.position_0_29\: out    vl_logic;
        \ball_next.position_0_30\: out    vl_logic;
        \ball_next.position_0_31\: out    vl_logic;
        \ball_next.radius\: out    vl_logic_vector(31 downto 0)
    );
end ball_move_computation;
